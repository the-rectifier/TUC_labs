LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY CLA_FA_TB IS
END CLA_FA_TB;
 
ARCHITECTURE behavior OF CLA_FA_TB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT CLA_FA
    PORT(
         A : IN  std_logic_vector(3 downto 0);
         B : IN  std_logic_vector(3 downto 0);
         Cin : IN  std_logic;
         S : OUT  std_logic_vector(3 downto 0);
		 Cout : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal A : std_logic_vector(3 downto 0) := (others => '0');
   signal B : std_logic_vector(3 downto 0) := (others => '0');
   signal Cin : std_logic := '0';

 	--Outputs
   signal Cout : std_logic;
   signal S : std_logic_vector(3 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: CLA_FA PORT MAP (
          A => A,
          B => B,
          Cin => Cin,
          S => S,
		  Cout => Cout
        );

   -- Clock process definitions


   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.

A <= X"0";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"0";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"0";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"1";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"1";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"2";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"2";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"3";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"3";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"4";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"4";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"5";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"5";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"6";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"6";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"7";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"7";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"8";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"8";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"9";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"9";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"a";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"a";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"b";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"b";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"c";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"c";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"d";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"d";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"e";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"e";
B <= X"f";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"0";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"0";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"1";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"1";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"2";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"2";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"3";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"3";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"4";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"4";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"5";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"5";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"6";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"6";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"7";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"7";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"8";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"8";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"9";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"9";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"a";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"a";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"b";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"b";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"c";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"c";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"d";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"d";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"e";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"e";
Cin <= '1';
wait for 1 ns;
A <= X"f";
B <= X"f";
Cin <= '0';
wait for 1 ns;
A <= X"f";
B <= X"f";
Cin <= '1';
wait for 1 ns;

      wait;
   end process;

END;
